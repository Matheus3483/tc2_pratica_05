`ifndef CDPRAM_SV
`define CDPRAM_SV


`define CDPRAM_SEL_CONTROL  0
`define CDPRAM_SEL_DATA_IN  1
`define CDPRAM_SEL_DATA_OUT 2
`define CDPRAM_SEL_STATUS   3


`endif